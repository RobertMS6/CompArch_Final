module processor()

endmodule